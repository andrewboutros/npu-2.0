module dsp_block_int8 # (
	parameter USE_CHAINADDER = "true",
	parameter IDATAW = 8,
	parameter ODATAW = 18
)(
	input clk,
	input rst,
	input [IDATAW-1:0] ax,
	input [IDATAW-1:0] ay,
	input [IDATAW-1:0] bx,
	input [IDATAW-1:0] by,
	input [IDATAW-1:0] cx,
	input [IDATAW-1:0] cy,
	input [IDATAW-1:0] dx,
	input [IDATAW-1:0] dy,
	input [63:0] chainin,
	output [63:0] chainout,
	output [ODATAW-1:0] resulta
);

tennm_mac tennm_mac_component (
	.ax (ax),
	.ay (ay),
	.bx (bx),
	.by (by),
	.chainin (chainin),
	.clr ({1'b0, 1'b0}),
	.clk (clk),
	.cx (cx),
	.cy (cy),
	.dx (dx),
	.dy (dy),
	.ena ({~rst, ~rst, ~rst}),
	.chainout (chainout),
	.resulta (resulta)
);

defparam
	tennm_mac_component.operation_mode = "m9x9_sumof4",
	tennm_mac_component.signed_max = "true",
	tennm_mac_component.signed_may = "true",
	tennm_mac_component.signed_mbx = "true",
	tennm_mac_component.signed_mby = "true",
	tennm_mac_component.signed_mcx = "true",
	tennm_mac_component.signed_mcy = "true",
	tennm_mac_component.signed_mdx = "true",
	tennm_mac_component.signed_mdy = "true",
	tennm_mac_component.sub_clken = "no_reg",
	tennm_mac_component.ay_use_scan_in = "false",
	tennm_mac_component.by_use_scan_in = "false",
	tennm_mac_component.delay_scan_out_ay = "false",
	tennm_mac_component.delay_scan_out_by = "false",
	tennm_mac_component.ax_width = IDATAW,
	tennm_mac_component.ax_clken = "0",
	tennm_mac_component.bx_width = IDATAW,
	tennm_mac_component.bx_clken = "0",
	tennm_mac_component.cx_width = IDATAW,
	tennm_mac_component.cx_clken = "0",
	tennm_mac_component.dx_width = IDATAW,
	tennm_mac_component.dx_clken = "0",
	tennm_mac_component.ay_scan_in_width = IDATAW,
	tennm_mac_component.ay_scan_in_clken = "0",
	tennm_mac_component.by_width = IDATAW,
	tennm_mac_component.by_clken = "0",
	tennm_mac_component.cy_width = IDATAW,
	tennm_mac_component.cy_clken = "0",
	tennm_mac_component.dy_width = IDATAW,
	tennm_mac_component.dy_clken = "0",
	tennm_mac_component.result_a_width = ODATAW,
	tennm_mac_component.output_clken = "0",
	tennm_mac_component.input_systolic_clken = "no_reg",
	tennm_mac_component.operand_source_may = "input",
	tennm_mac_component.operand_source_mby = "input",
	tennm_mac_component.preadder_subtract_a = "false",
	tennm_mac_component.preadder_subtract_b = "false",
	tennm_mac_component.az_clken = "no_reg",
	tennm_mac_component.bz_clken = "no_reg",
	tennm_mac_component.operand_source_max = "input",
	tennm_mac_component.operand_source_mbx = "input",
	tennm_mac_component.coef_sel_a_clken = "no_reg",
	tennm_mac_component.coef_sel_b_clken = "no_reg",
	tennm_mac_component.coef_a_0 = 0,
	tennm_mac_component.coef_a_1 = 0,
	tennm_mac_component.coef_a_2 = 0,
	tennm_mac_component.coef_a_3 = 0,
	tennm_mac_component.coef_a_4 = 0,
	tennm_mac_component.coef_a_5 = 0,
	tennm_mac_component.coef_a_6 = 0,
	tennm_mac_component.coef_a_7 = 0,
	tennm_mac_component.coef_b_0 = 0,
	tennm_mac_component.coef_b_1 = 0,
	tennm_mac_component.coef_b_2 = 0,
	tennm_mac_component.coef_b_3 = 0,
	tennm_mac_component.coef_b_4 = 0,
	tennm_mac_component.coef_b_5 = 0,
	tennm_mac_component.coef_b_6 = 0,
	tennm_mac_component.coef_b_7 = 0,
	tennm_mac_component.accumulate_clken = "no_reg",
	tennm_mac_component.load_const_clken = "no_reg",
	tennm_mac_component.negate_clken = "no_reg",
	tennm_mac_component.enable_double_accum = "false",
	tennm_mac_component.load_const_value = 0,
	tennm_mac_component.use_chainadder = USE_CHAINADDER,
	tennm_mac_component.chain_inout_width = 64,
	tennm_mac_component.input_pipeline_clken = "0",
	tennm_mac_component.second_pipeline_clken = "0",
	tennm_mac_component.accum_pipeline_clken = "no_reg",
	tennm_mac_component.accum_2nd_pipeline_clken = "no_reg",
	tennm_mac_component.load_const_pipeline_clken = "no_reg",
	tennm_mac_component.load_const_2nd_pipeline_clken = "no_reg",
	tennm_mac_component.clear_type = "none";
			  
endmodule